-- sopc_compteur
