-- sopc_compteur